module fx_to_ft
  (
    input logic [23:0] x,
    output logic [31:0] y
  );

  logic [22:0] no_sign;
  logic [22:0] mantissa;
  logic [7:0] exponent;

  int unsigned leading_zeros;

  always_comb begin
    no_sign = 23'(x[23] ? ~x[22:0] + 1 : x[22:0]);
    leading_zeros = 0;

  // DOES NOT MEET TIMING

    // if (no_sign != 23'b0) begin
    //   for (int i = 0; i < 22; i++) begin
    //     if (no_sign[22 - i] == 1'b1) begin
    //       break;
    //     end
    //     else begin
    //       leading_zeros++;
    //     end
    //   end
    // end

    // leading_zeros = no_sign[22] ? 0 : no_sign[21] ? 1 : 2;

    casex(no_sign) 
      23'b00000000000000000000001: leading_zeros = 22;
      23'b0000000000000000000001?: leading_zeros = 21;
      23'b000000000000000000001??: leading_zeros = 20;
      23'b00000000000000000001???: leading_zeros = 19;
      23'b0000000000000000001????: leading_zeros = 18;
      23'b000000000000000001?????: leading_zeros = 17;
      23'b00000000000000001??????: leading_zeros = 16;
      23'b0000000000000001???????: leading_zeros = 15;
      23'b000000000000001????????: leading_zeros = 14;
      23'b00000000000001?????????: leading_zeros = 13;
      23'b0000000000001??????????: leading_zeros = 12;
      23'b000000000001???????????: leading_zeros = 11;
      23'b00000000001????????????: leading_zeros = 10;
      23'b0000000001?????????????: leading_zeros = 9;
      23'b000000001??????????????: leading_zeros = 8;
      23'b00000001???????????????: leading_zeros = 7;
      23'b0000001????????????????: leading_zeros = 6;
      23'b000001?????????????????: leading_zeros = 5;
      23'b00001??????????????????: leading_zeros = 4;
      23'b0001???????????????????: leading_zeros = 3;
      23'b001????????????????????: leading_zeros = 2;
      23'b01?????????????????????: leading_zeros = 1;
      default: leading_zeros = 0;
    endcase

    mantissa = no_sign << (leading_zeros + 1); // exclude MSB

    exponent = 8'(127 - leading_zeros);

    y = {x[23], exponent, mantissa};
  end
endmodule